.title KiCad schematic
V1 Net-_V1-Pad1_ 0 dc(12)
V2 E22-PG 0 pulse(0 3 2n 2n 2n 60ms 180ms)
V4 E21-PG 0 pulse(0 3 90ms 2n 2n 60ms 180ms)
VBOGUS1 Net-_V1-Pad1_ E24-12V dc(0)
R1 Net-_D1-Pad1_ E22-PG 3k
Q1 FF1 Net-_D1-Pad2_ 0 BCY58
R2 FF2 E22-PG 3k
D1 Net-_D1-Pad1_ Net-_D1-Pad2_ DIODE
R5 Net-_C1-Pad1_ Net-_D1-Pad2_ 300
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 2n2
D2 Net-_D2-Pad1_ Net-_C1-Pad2_ DIODE
R4 Net-_D2-Pad1_ E21-PG 3k
R3 FF1 E21-PG 3k
R6 0 Net-_D1-Pad2_ 180k
R8 FF1 E24-12V 1k
Q2 FF2 Net-_C1-Pad2_ 0 BCY58
R7 0 Net-_C1-Pad2_ 180k
R9 FF2 E24-12V 1k
R10 Net-_Q3-Pad2_ FF1 10k
Q3 Net-_Q3-Pad1_ Net-_Q3-Pad2_ 0 BCY58
R12 Net-_Q3-Pad1_ E24-12V 2k
R13 INT-7 Net-_Q3-Pad1_ 5k1
R15 INT-7 Net-_Q4-Pad1_ 5k1
R14 Net-_Q4-Pad1_ E24-12V 2k
Q4 Net-_Q4-Pad1_ Net-_Q4-Pad2_ 0 BCY58
R11 Net-_Q4-Pad2_ FF2 10k
R16 Net-_D3-Pad1_ E14-PG 3k
Q5 FF3 Net-_D3-Pad2_ 0 BCY58
R17 FF4 E14-PG 3k
D3 Net-_D3-Pad1_ Net-_D3-Pad2_ DIODE
R20 Net-_C2-Pad1_ Net-_D3-Pad2_ 300
C2 Net-_C2-Pad1_ Net-_C2-Pad2_ 2n2
D4 Net-_D4-Pad1_ Net-_C2-Pad2_ DIODE
R19 Net-_D4-Pad1_ E13-PG 3k
R18 FF3 E13-PG 3k
R21 0 Net-_D3-Pad2_ 180k
R23 FF3 E24-12V 1k
Q6 FF4 Net-_C2-Pad2_ 0 BCY58
R22 0 Net-_C2-Pad2_ 180k
R24 FF4 E24-12V 1k
R25 Net-_Q4-Pad2_ FF3 10k
R26 Net-_Q3-Pad2_ FF4 10k
V3 E14-PG 0 pulse(0 3 45ms 2n 2n 60ms 180ms)
V5 E13-PG 0 pulse(0 3 135ms 2n 2n 60ms 180ms)
R27 AUX12-TGL E24-12V 1k
Q7 AUX12-TGL INT-7 0 BCY58
Q8 AUX11-TGL Net-_Q8-Pad2_ 0 BCY58
R28 Net-_Q8-Pad2_ AUX12-TGL 10k
R29 AUX11-TGL E24-12V 1k
.model DIODE D 
.model BCY58 npn 
.model BSX95 npn 
.model AUY21 pnp 
.tran 1ms 600ms 120m 
.control 
run 
rusage 
set filetype=ascii 
set color0=white 
set xbrushwidth=5 
write "C:\Users\andy\OneDrive\Documents\MPS Tune-o-Matic\trunk\Simulation\Pressure Loop\PressureLoop.out" "V(E22-PG)" "V(E21-PG)" "V(E14-PG)" "V(E13-PG)" "V(INT-7)" 
plot "V(E22-PG)"+5 "V(E14-PG)"+10 "V(E21-PG)"+15 "V(E13-PG)"+20 "V(INT-7)" 
.endc 
.end
