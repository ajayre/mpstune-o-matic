.title KiCad schematic
.include "MPS.lib"
V2 Net-_V2-Pad1_ 0 dc(12)
VBOGUS2 Net-_V2-Pad1_ E24-12V dc(0)
R48 AUX12-TGL E24-12V 1k
Q8 AUX12-TGL IN 0 BCY58
Q10 AUX11-TGL Net-_Q10-Pad2_ 0 BCY58
R50 Net-_Q10-Pad2_ AUX12-TGL 10k
R53 AUX11-TGL E24-12V 1k
C5 AUX11-TGL Net-_C5-Pad2_ 6.8n
R30 Net-_C4-Pad2_ AUX1-10V 130k
R31 0 Net-_C4-Pad2_ 68k
D4 EDGES Net-_C4-Pad2_ DIODE
R26 0 Net-_C5-Pad2_ 68k
R25 Net-_C5-Pad2_ AUX1-10V 130k
D5 EDGES Net-_C5-Pad2_ DIODE
R23 EDGES AUX1-10V 100k
VBOGUS1 Net-_V1-Pad1_ AUX1-10V dc(0)
V1 Net-_V1-Pad1_ 0 dc(10)
D15 EDGES E8-MPS DIODE
D16 EDGES Net-_D16-Pad2_ DIODE
Q11 AUX10-SP Net-_D16-Pad2_ 0 BCY58
R65 0 Net-_D16-Pad2_ 180k
R68 Net-_C9-Pad2_ Net-_D16-Pad2_ 300
C9 Net-_C9-Pad1_ Net-_C9-Pad2_ 1.0n
R67 Net-_C9-Pad1_ AUX10-SP 2k4
Q12 BASE_PULSE Net-_C9-Pad1_ 0 BCY58
R66 AUX10-SP AUX1-10V 2k
R69 BASE_PULSE AUX1-10V 1k
R64 E15-MPS AUX1-10V 510
R63 E15-MPS Net-_D14-Pad2_ 2k2
D14 Net-_D14-Pad1_ Net-_D14-Pad2_ DIODE
R62 Net-_D14-Pad1_ AUX1-10V 1k2
R61 Net-_D14-Pad1_ E1-T1 240
V7 INT-6 0 dc(5.0)
XTR1 BASE_PULSE E15-MPS E8-MPS E10-MPS mps vac=15
C4 AUX12-TGL Net-_C4-Pad2_ 6.8n
V8 IN 0 pulse(0 5 2n 2n 2n 3ms 6ms)
Q1 Net-_Q1-Pad1_ Net-_Q1-Pad2_ 0 BCY58
R2 BASE_PULSE Net-_Q1-Pad2_ 20k
R1 Net-_Q1-Pad1_ AUX1-10V 2k
R3 Net-_Q1-Pad2_ 0 10k
R4 OUT Net-_Q1-Pad1_ 10k
R5 0 OUT 12k
R7 0 E10-MPS 1k
RV1 INT-6 E10-MPS 5k
RV2 E1-T1 0 1k
.model DIODE D 
.model BCY58 npn 
.model BSX95 npn 
.model AUY21 pnp 
.tran 0.05ms 100ms 89m 
.control 
run 
rusage 
set filetype=ascii 
set color0=white 
set xbrushwidth=5 
*write "C:\Users\andy\OneDrive\Documents\MPS Tune-o-Matic\trunk\Simulation\Pressure Loop\PressureLoop.out" "V(BASE_PULSE)" "V(INT-7)" 
plot "V(IN)"+0 "V(BASE_PULSE)"+6 "V(OUT)"+33 
.endc 
.end
